VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO R4_butter
  CLASS BLOCK ;
  FOREIGN R4_butter ;
  ORIGIN 0.000 0.000 ;
  SIZE 300.000 BY 200.000 ;
  PIN Xio[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 49.680 300.000 50.280 ;
    END
  END Xio[0]
  PIN Xio[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 97.280 300.000 97.880 ;
    END
  END Xio[1]
  PIN Xio[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 144.880 300.000 145.480 ;
    END
  END Xio[2]
  PIN Xio[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 192.480 300.000 193.080 ;
    END
  END Xio[3]
  PIN Xro[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 44.920 300.000 45.520 ;
    END
  END Xro[0]
  PIN Xro[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 92.520 300.000 93.120 ;
    END
  END Xro[1]
  PIN Xro[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 140.120 300.000 140.720 ;
    END
  END Xro[2]
  PIN Xro[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 187.720 300.000 188.320 ;
    END
  END Xro[3]
  PIN c1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 165.960 4.000 166.560 ;
    END
  END c1
  PIN c2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 99.320 4.000 99.920 ;
    END
  END c2
  PIN c3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 32.680 4.000 33.280 ;
    END
  END c3
  PIN la_oenb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 37.350 0.000 37.630 4.000 ;
    END
  END la_oenb[0]
  PIN la_oenb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 112.330 0.000 112.610 4.000 ;
    END
  END la_oenb[1]
  PIN la_oenb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 187.310 0.000 187.590 4.000 ;
    END
  END la_oenb[2]
  PIN la_oenb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 262.290 0.000 262.570 4.000 ;
    END
  END la_oenb[3]
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 187.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 187.920 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 187.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 187.920 ;
    END
  END vssd1
  PIN xi0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 11.600 300.000 12.200 ;
    END
  END xi0[0]
  PIN xi0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 59.200 300.000 59.800 ;
    END
  END xi0[1]
  PIN xi0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 106.800 300.000 107.400 ;
    END
  END xi0[2]
  PIN xi0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 154.400 300.000 155.000 ;
    END
  END xi0[3]
  PIN xi1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 21.120 300.000 21.720 ;
    END
  END xi1[0]
  PIN xi1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 68.720 300.000 69.320 ;
    END
  END xi1[1]
  PIN xi1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 116.320 300.000 116.920 ;
    END
  END xi1[2]
  PIN xi1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 163.920 300.000 164.520 ;
    END
  END xi1[3]
  PIN xi2[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 30.640 300.000 31.240 ;
    END
  END xi2[0]
  PIN xi2[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 78.240 300.000 78.840 ;
    END
  END xi2[1]
  PIN xi2[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 125.840 300.000 126.440 ;
    END
  END xi2[2]
  PIN xi2[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 173.440 300.000 174.040 ;
    END
  END xi2[3]
  PIN xi3[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 40.160 300.000 40.760 ;
    END
  END xi3[0]
  PIN xi3[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 87.760 300.000 88.360 ;
    END
  END xi3[1]
  PIN xi3[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 135.360 300.000 135.960 ;
    END
  END xi3[2]
  PIN xi3[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 182.960 300.000 183.560 ;
    END
  END xi3[3]
  PIN xr0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 6.840 300.000 7.440 ;
    END
  END xr0[0]
  PIN xr0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 54.440 300.000 55.040 ;
    END
  END xr0[1]
  PIN xr0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 102.040 300.000 102.640 ;
    END
  END xr0[2]
  PIN xr0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 149.640 300.000 150.240 ;
    END
  END xr0[3]
  PIN xr1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 16.360 300.000 16.960 ;
    END
  END xr1[0]
  PIN xr1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 63.960 300.000 64.560 ;
    END
  END xr1[1]
  PIN xr1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 111.560 300.000 112.160 ;
    END
  END xr1[2]
  PIN xr1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 159.160 300.000 159.760 ;
    END
  END xr1[3]
  PIN xr2[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 25.880 300.000 26.480 ;
    END
  END xr2[0]
  PIN xr2[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 73.480 300.000 74.080 ;
    END
  END xr2[1]
  PIN xr2[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 121.080 300.000 121.680 ;
    END
  END xr2[2]
  PIN xr2[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 168.680 300.000 169.280 ;
    END
  END xr2[3]
  PIN xr3[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 35.400 300.000 36.000 ;
    END
  END xr3[0]
  PIN xr3[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 83.000 300.000 83.600 ;
    END
  END xr3[1]
  PIN xr3[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 130.600 300.000 131.200 ;
    END
  END xr3[2]
  PIN xr3[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 178.200 300.000 178.800 ;
    END
  END xr3[3]
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 294.400 187.765 ;
      LAYER met1 ;
        RECT 4.670 10.640 295.250 187.920 ;
      LAYER met2 ;
        RECT 4.690 4.280 295.230 192.965 ;
        RECT 4.690 4.000 37.070 4.280 ;
        RECT 37.910 4.000 112.050 4.280 ;
        RECT 112.890 4.000 187.030 4.280 ;
        RECT 187.870 4.000 262.010 4.280 ;
        RECT 262.850 4.000 295.230 4.280 ;
      LAYER met3 ;
        RECT 4.000 192.080 295.600 192.945 ;
        RECT 4.000 188.720 296.000 192.080 ;
        RECT 4.000 187.320 295.600 188.720 ;
        RECT 4.000 183.960 296.000 187.320 ;
        RECT 4.000 182.560 295.600 183.960 ;
        RECT 4.000 179.200 296.000 182.560 ;
        RECT 4.000 177.800 295.600 179.200 ;
        RECT 4.000 174.440 296.000 177.800 ;
        RECT 4.000 173.040 295.600 174.440 ;
        RECT 4.000 169.680 296.000 173.040 ;
        RECT 4.000 168.280 295.600 169.680 ;
        RECT 4.000 166.960 296.000 168.280 ;
        RECT 4.400 165.560 296.000 166.960 ;
        RECT 4.000 164.920 296.000 165.560 ;
        RECT 4.000 163.520 295.600 164.920 ;
        RECT 4.000 160.160 296.000 163.520 ;
        RECT 4.000 158.760 295.600 160.160 ;
        RECT 4.000 155.400 296.000 158.760 ;
        RECT 4.000 154.000 295.600 155.400 ;
        RECT 4.000 150.640 296.000 154.000 ;
        RECT 4.000 149.240 295.600 150.640 ;
        RECT 4.000 145.880 296.000 149.240 ;
        RECT 4.000 144.480 295.600 145.880 ;
        RECT 4.000 141.120 296.000 144.480 ;
        RECT 4.000 139.720 295.600 141.120 ;
        RECT 4.000 136.360 296.000 139.720 ;
        RECT 4.000 134.960 295.600 136.360 ;
        RECT 4.000 131.600 296.000 134.960 ;
        RECT 4.000 130.200 295.600 131.600 ;
        RECT 4.000 126.840 296.000 130.200 ;
        RECT 4.000 125.440 295.600 126.840 ;
        RECT 4.000 122.080 296.000 125.440 ;
        RECT 4.000 120.680 295.600 122.080 ;
        RECT 4.000 117.320 296.000 120.680 ;
        RECT 4.000 115.920 295.600 117.320 ;
        RECT 4.000 112.560 296.000 115.920 ;
        RECT 4.000 111.160 295.600 112.560 ;
        RECT 4.000 107.800 296.000 111.160 ;
        RECT 4.000 106.400 295.600 107.800 ;
        RECT 4.000 103.040 296.000 106.400 ;
        RECT 4.000 101.640 295.600 103.040 ;
        RECT 4.000 100.320 296.000 101.640 ;
        RECT 4.400 98.920 296.000 100.320 ;
        RECT 4.000 98.280 296.000 98.920 ;
        RECT 4.000 96.880 295.600 98.280 ;
        RECT 4.000 93.520 296.000 96.880 ;
        RECT 4.000 92.120 295.600 93.520 ;
        RECT 4.000 88.760 296.000 92.120 ;
        RECT 4.000 87.360 295.600 88.760 ;
        RECT 4.000 84.000 296.000 87.360 ;
        RECT 4.000 82.600 295.600 84.000 ;
        RECT 4.000 79.240 296.000 82.600 ;
        RECT 4.000 77.840 295.600 79.240 ;
        RECT 4.000 74.480 296.000 77.840 ;
        RECT 4.000 73.080 295.600 74.480 ;
        RECT 4.000 69.720 296.000 73.080 ;
        RECT 4.000 68.320 295.600 69.720 ;
        RECT 4.000 64.960 296.000 68.320 ;
        RECT 4.000 63.560 295.600 64.960 ;
        RECT 4.000 60.200 296.000 63.560 ;
        RECT 4.000 58.800 295.600 60.200 ;
        RECT 4.000 55.440 296.000 58.800 ;
        RECT 4.000 54.040 295.600 55.440 ;
        RECT 4.000 50.680 296.000 54.040 ;
        RECT 4.000 49.280 295.600 50.680 ;
        RECT 4.000 45.920 296.000 49.280 ;
        RECT 4.000 44.520 295.600 45.920 ;
        RECT 4.000 41.160 296.000 44.520 ;
        RECT 4.000 39.760 295.600 41.160 ;
        RECT 4.000 36.400 296.000 39.760 ;
        RECT 4.000 35.000 295.600 36.400 ;
        RECT 4.000 33.680 296.000 35.000 ;
        RECT 4.400 32.280 296.000 33.680 ;
        RECT 4.000 31.640 296.000 32.280 ;
        RECT 4.000 30.240 295.600 31.640 ;
        RECT 4.000 26.880 296.000 30.240 ;
        RECT 4.000 25.480 295.600 26.880 ;
        RECT 4.000 22.120 296.000 25.480 ;
        RECT 4.000 20.720 295.600 22.120 ;
        RECT 4.000 17.360 296.000 20.720 ;
        RECT 4.000 15.960 295.600 17.360 ;
        RECT 4.000 12.600 296.000 15.960 ;
        RECT 4.000 11.200 295.600 12.600 ;
        RECT 4.000 7.840 296.000 11.200 ;
        RECT 4.000 6.975 295.600 7.840 ;
  END
END R4_butter
END LIBRARY

