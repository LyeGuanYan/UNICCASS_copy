magic
tech sky130A
magscale 1 2
timestamp 1697601861
<< obsli1 >>
rect 1104 2159 35236 36465
<< obsm1 >>
rect 934 2128 35590 36496
<< metal2 >>
rect 4526 0 4582 800
rect 13634 0 13690 800
rect 22742 0 22798 800
rect 31850 0 31906 800
<< obsm2 >>
rect 938 856 35584 37913
rect 938 711 4470 856
rect 4638 711 13578 856
rect 13746 711 22686 856
rect 22854 711 31794 856
rect 31962 711 35584 856
<< metal3 >>
rect 35600 37816 36400 37936
rect 35600 36864 36400 36984
rect 35600 35912 36400 36032
rect 35600 34960 36400 35080
rect 35600 34008 36400 34128
rect 35600 33056 36400 33176
rect 0 32240 800 32360
rect 35600 32104 36400 32224
rect 35600 31152 36400 31272
rect 35600 30200 36400 30320
rect 35600 29248 36400 29368
rect 35600 28296 36400 28416
rect 35600 27344 36400 27464
rect 35600 26392 36400 26512
rect 35600 25440 36400 25560
rect 35600 24488 36400 24608
rect 35600 23536 36400 23656
rect 35600 22584 36400 22704
rect 35600 21632 36400 21752
rect 35600 20680 36400 20800
rect 35600 19728 36400 19848
rect 0 19320 800 19440
rect 35600 18776 36400 18896
rect 35600 17824 36400 17944
rect 35600 16872 36400 16992
rect 35600 15920 36400 16040
rect 35600 14968 36400 15088
rect 35600 14016 36400 14136
rect 35600 13064 36400 13184
rect 35600 12112 36400 12232
rect 35600 11160 36400 11280
rect 35600 10208 36400 10328
rect 35600 9256 36400 9376
rect 35600 8304 36400 8424
rect 35600 7352 36400 7472
rect 0 6400 800 6520
rect 35600 6400 36400 6520
rect 35600 5448 36400 5568
rect 35600 4496 36400 4616
rect 35600 3544 36400 3664
rect 35600 2592 36400 2712
rect 35600 1640 36400 1760
rect 35600 688 36400 808
<< obsm3 >>
rect 800 37736 35520 37909
rect 800 37064 35600 37736
rect 800 36784 35520 37064
rect 800 36112 35600 36784
rect 800 35832 35520 36112
rect 800 35160 35600 35832
rect 800 34880 35520 35160
rect 800 34208 35600 34880
rect 800 33928 35520 34208
rect 800 33256 35600 33928
rect 800 32976 35520 33256
rect 800 32440 35600 32976
rect 880 32304 35600 32440
rect 880 32160 35520 32304
rect 800 32024 35520 32160
rect 800 31352 35600 32024
rect 800 31072 35520 31352
rect 800 30400 35600 31072
rect 800 30120 35520 30400
rect 800 29448 35600 30120
rect 800 29168 35520 29448
rect 800 28496 35600 29168
rect 800 28216 35520 28496
rect 800 27544 35600 28216
rect 800 27264 35520 27544
rect 800 26592 35600 27264
rect 800 26312 35520 26592
rect 800 25640 35600 26312
rect 800 25360 35520 25640
rect 800 24688 35600 25360
rect 800 24408 35520 24688
rect 800 23736 35600 24408
rect 800 23456 35520 23736
rect 800 22784 35600 23456
rect 800 22504 35520 22784
rect 800 21832 35600 22504
rect 800 21552 35520 21832
rect 800 20880 35600 21552
rect 800 20600 35520 20880
rect 800 19928 35600 20600
rect 800 19648 35520 19928
rect 800 19520 35600 19648
rect 880 19240 35600 19520
rect 800 18976 35600 19240
rect 800 18696 35520 18976
rect 800 18024 35600 18696
rect 800 17744 35520 18024
rect 800 17072 35600 17744
rect 800 16792 35520 17072
rect 800 16120 35600 16792
rect 800 15840 35520 16120
rect 800 15168 35600 15840
rect 800 14888 35520 15168
rect 800 14216 35600 14888
rect 800 13936 35520 14216
rect 800 13264 35600 13936
rect 800 12984 35520 13264
rect 800 12312 35600 12984
rect 800 12032 35520 12312
rect 800 11360 35600 12032
rect 800 11080 35520 11360
rect 800 10408 35600 11080
rect 800 10128 35520 10408
rect 800 9456 35600 10128
rect 800 9176 35520 9456
rect 800 8504 35600 9176
rect 800 8224 35520 8504
rect 800 7552 35600 8224
rect 800 7272 35520 7552
rect 800 6600 35600 7272
rect 880 6320 35520 6600
rect 800 5648 35600 6320
rect 800 5368 35520 5648
rect 800 4696 35600 5368
rect 800 4416 35520 4696
rect 800 3744 35600 4416
rect 800 3464 35520 3744
rect 800 2792 35600 3464
rect 800 2512 35520 2792
rect 800 1840 35600 2512
rect 800 1560 35520 1840
rect 800 888 35600 1560
rect 800 715 35520 888
<< metal4 >>
rect 4208 2128 4528 36496
rect 19568 2128 19888 36496
rect 34928 2128 35248 36496
<< labels >>
rlabel metal3 s 35600 9256 36400 9376 6 Xio[0]
port 1 nsew signal output
rlabel metal3 s 35600 18776 36400 18896 6 Xio[1]
port 2 nsew signal output
rlabel metal3 s 35600 28296 36400 28416 6 Xio[2]
port 3 nsew signal output
rlabel metal3 s 35600 37816 36400 37936 6 Xio[3]
port 4 nsew signal output
rlabel metal3 s 35600 8304 36400 8424 6 Xro[0]
port 5 nsew signal output
rlabel metal3 s 35600 17824 36400 17944 6 Xro[1]
port 6 nsew signal output
rlabel metal3 s 35600 27344 36400 27464 6 Xro[2]
port 7 nsew signal output
rlabel metal3 s 35600 36864 36400 36984 6 Xro[3]
port 8 nsew signal output
rlabel metal3 s 0 32240 800 32360 6 c1
port 9 nsew signal input
rlabel metal3 s 0 19320 800 19440 6 c2
port 10 nsew signal input
rlabel metal3 s 0 6400 800 6520 6 c3
port 11 nsew signal input
rlabel metal2 s 4526 0 4582 800 6 la_oenb[0]
port 12 nsew signal output
rlabel metal2 s 13634 0 13690 800 6 la_oenb[1]
port 13 nsew signal output
rlabel metal2 s 22742 0 22798 800 6 la_oenb[2]
port 14 nsew signal output
rlabel metal2 s 31850 0 31906 800 6 la_oenb[3]
port 15 nsew signal output
rlabel metal4 s 4208 2128 4528 36496 6 vccd1
port 16 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 36496 6 vccd1
port 16 nsew power bidirectional
rlabel metal4 s 19568 2128 19888 36496 6 vssd1
port 17 nsew ground bidirectional
rlabel metal3 s 35600 1640 36400 1760 6 xi0[0]
port 18 nsew signal input
rlabel metal3 s 35600 11160 36400 11280 6 xi0[1]
port 19 nsew signal input
rlabel metal3 s 35600 20680 36400 20800 6 xi0[2]
port 20 nsew signal input
rlabel metal3 s 35600 30200 36400 30320 6 xi0[3]
port 21 nsew signal input
rlabel metal3 s 35600 3544 36400 3664 6 xi1[0]
port 22 nsew signal input
rlabel metal3 s 35600 13064 36400 13184 6 xi1[1]
port 23 nsew signal input
rlabel metal3 s 35600 22584 36400 22704 6 xi1[2]
port 24 nsew signal input
rlabel metal3 s 35600 32104 36400 32224 6 xi1[3]
port 25 nsew signal input
rlabel metal3 s 35600 5448 36400 5568 6 xi2[0]
port 26 nsew signal input
rlabel metal3 s 35600 14968 36400 15088 6 xi2[1]
port 27 nsew signal input
rlabel metal3 s 35600 24488 36400 24608 6 xi2[2]
port 28 nsew signal input
rlabel metal3 s 35600 34008 36400 34128 6 xi2[3]
port 29 nsew signal input
rlabel metal3 s 35600 7352 36400 7472 6 xi3[0]
port 30 nsew signal input
rlabel metal3 s 35600 16872 36400 16992 6 xi3[1]
port 31 nsew signal input
rlabel metal3 s 35600 26392 36400 26512 6 xi3[2]
port 32 nsew signal input
rlabel metal3 s 35600 35912 36400 36032 6 xi3[3]
port 33 nsew signal input
rlabel metal3 s 35600 688 36400 808 6 xr0[0]
port 34 nsew signal input
rlabel metal3 s 35600 10208 36400 10328 6 xr0[1]
port 35 nsew signal input
rlabel metal3 s 35600 19728 36400 19848 6 xr0[2]
port 36 nsew signal input
rlabel metal3 s 35600 29248 36400 29368 6 xr0[3]
port 37 nsew signal input
rlabel metal3 s 35600 2592 36400 2712 6 xr1[0]
port 38 nsew signal input
rlabel metal3 s 35600 12112 36400 12232 6 xr1[1]
port 39 nsew signal input
rlabel metal3 s 35600 21632 36400 21752 6 xr1[2]
port 40 nsew signal input
rlabel metal3 s 35600 31152 36400 31272 6 xr1[3]
port 41 nsew signal input
rlabel metal3 s 35600 4496 36400 4616 6 xr2[0]
port 42 nsew signal input
rlabel metal3 s 35600 14016 36400 14136 6 xr2[1]
port 43 nsew signal input
rlabel metal3 s 35600 23536 36400 23656 6 xr2[2]
port 44 nsew signal input
rlabel metal3 s 35600 33056 36400 33176 6 xr2[3]
port 45 nsew signal input
rlabel metal3 s 35600 6400 36400 6520 6 xr3[0]
port 46 nsew signal input
rlabel metal3 s 35600 15920 36400 16040 6 xr3[1]
port 47 nsew signal input
rlabel metal3 s 35600 25440 36400 25560 6 xr3[2]
port 48 nsew signal input
rlabel metal3 s 35600 34960 36400 35080 6 xr3[3]
port 49 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 36400 38800
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 445408
string GDS_FILE /home/guanyanlye/unic-cass/caravel_tutorial/caravel_uniccas_example/openlane/R4_butter/runs/23_10_18_12_03/results/signoff/R4_butter.magic.gds
string GDS_START 56748
<< end >>

