magic
tech sky130A
magscale 1 2
timestamp 1699459426
<< nwell >>
rect 1066 36165 35274 36486
rect 1066 35077 35274 35643
rect 1066 33989 35274 34555
rect 1066 32901 35274 33467
rect 1066 31813 35274 32379
rect 1066 30725 35274 31291
rect 1066 29637 35274 30203
rect 1066 28549 35274 29115
rect 1066 27461 35274 28027
rect 1066 26373 35274 26939
rect 1066 25285 35274 25851
rect 1066 24197 35274 24763
rect 1066 23109 35274 23675
rect 1066 22021 35274 22587
rect 1066 20933 35274 21499
rect 1066 19845 35274 20411
rect 1066 18757 35274 19323
rect 1066 17669 35274 18235
rect 1066 16581 35274 17147
rect 1066 15493 35274 16059
rect 1066 14405 35274 14971
rect 1066 13317 35274 13883
rect 1066 12229 35274 12795
rect 1066 11141 35274 11707
rect 1066 10053 35274 10619
rect 1066 8965 35274 9531
rect 1066 7877 35274 8443
rect 1066 6789 35274 7355
rect 1066 5701 35274 6267
rect 1066 4613 35274 5179
rect 1066 3525 35274 4091
rect 1066 2437 35274 3003
<< obsli1 >>
rect 1104 2159 35236 36465
<< obsm1 >>
rect 1104 76 35498 36496
<< metal2 >>
rect 1582 0 1638 800
rect 2410 0 2466 800
rect 3238 0 3294 800
rect 4066 0 4122 800
rect 4894 0 4950 800
rect 5722 0 5778 800
rect 6550 0 6606 800
rect 7378 0 7434 800
rect 8206 0 8262 800
rect 9034 0 9090 800
rect 9862 0 9918 800
rect 10690 0 10746 800
rect 11518 0 11574 800
rect 12346 0 12402 800
rect 13174 0 13230 800
rect 14002 0 14058 800
rect 14830 0 14886 800
rect 15658 0 15714 800
rect 16486 0 16542 800
rect 17314 0 17370 800
rect 18142 0 18198 800
rect 18970 0 19026 800
rect 19798 0 19854 800
rect 20626 0 20682 800
rect 21454 0 21510 800
rect 22282 0 22338 800
rect 23110 0 23166 800
rect 23938 0 23994 800
rect 24766 0 24822 800
rect 25594 0 25650 800
rect 26422 0 26478 800
rect 27250 0 27306 800
rect 28078 0 28134 800
rect 28906 0 28962 800
rect 29734 0 29790 800
rect 30562 0 30618 800
rect 31390 0 31446 800
rect 32218 0 32274 800
rect 33046 0 33102 800
rect 33874 0 33930 800
rect 34702 0 34758 800
<< obsm2 >>
rect 1584 856 35494 36485
rect 1694 70 2354 856
rect 2522 70 3182 856
rect 3350 70 4010 856
rect 4178 70 4838 856
rect 5006 70 5666 856
rect 5834 70 6494 856
rect 6662 70 7322 856
rect 7490 70 8150 856
rect 8318 70 8978 856
rect 9146 70 9806 856
rect 9974 70 10634 856
rect 10802 70 11462 856
rect 11630 70 12290 856
rect 12458 70 13118 856
rect 13286 70 13946 856
rect 14114 70 14774 856
rect 14942 70 15602 856
rect 15770 70 16430 856
rect 16598 70 17258 856
rect 17426 70 18086 856
rect 18254 70 18914 856
rect 19082 70 19742 856
rect 19910 70 20570 856
rect 20738 70 21398 856
rect 21566 70 22226 856
rect 22394 70 23054 856
rect 23222 70 23882 856
rect 24050 70 24710 856
rect 24878 70 25538 856
rect 25706 70 26366 856
rect 26534 70 27194 856
rect 27362 70 28022 856
rect 28190 70 28850 856
rect 29018 70 29678 856
rect 29846 70 30506 856
rect 30674 70 31334 856
rect 31502 70 32162 856
rect 32330 70 32990 856
rect 33158 70 33818 856
rect 33986 70 34646 856
rect 34814 70 35494 856
<< metal3 >>
rect 35600 33736 36400 33856
rect 35600 24080 36400 24200
rect 35600 14424 36400 14544
rect 35600 4768 36400 4888
<< obsm3 >>
rect 4210 33936 35600 36481
rect 4210 33656 35520 33936
rect 4210 24280 35600 33656
rect 4210 24000 35520 24280
rect 4210 14624 35600 24000
rect 4210 14344 35520 14624
rect 4210 4968 35600 14344
rect 4210 4688 35520 4968
rect 4210 2143 35600 4688
<< metal4 >>
rect 4208 2128 4528 36496
rect 19568 2128 19888 36496
rect 34928 2128 35248 36496
<< labels >>
rlabel metal2 s 34702 0 34758 800 6 CLK
port 1 nsew signal input
rlabel metal3 s 35600 33736 36400 33856 6 RST
port 2 nsew signal input
rlabel metal2 s 28906 0 28962 800 6 Xio[0]
port 3 nsew signal output
rlabel metal2 s 30562 0 30618 800 6 Xio[1]
port 4 nsew signal output
rlabel metal2 s 32218 0 32274 800 6 Xio[2]
port 5 nsew signal output
rlabel metal2 s 33874 0 33930 800 6 Xio[3]
port 6 nsew signal output
rlabel metal2 s 28078 0 28134 800 6 Xro[0]
port 7 nsew signal output
rlabel metal2 s 29734 0 29790 800 6 Xro[1]
port 8 nsew signal output
rlabel metal2 s 31390 0 31446 800 6 Xro[2]
port 9 nsew signal output
rlabel metal2 s 33046 0 33102 800 6 Xro[3]
port 10 nsew signal output
rlabel metal3 s 35600 4768 36400 4888 6 c1
port 11 nsew signal input
rlabel metal3 s 35600 14424 36400 14544 6 c2
port 12 nsew signal input
rlabel metal3 s 35600 24080 36400 24200 6 c3
port 13 nsew signal input
rlabel metal4 s 4208 2128 4528 36496 6 vccd1
port 14 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 36496 6 vccd1
port 14 nsew power bidirectional
rlabel metal4 s 19568 2128 19888 36496 6 vssd1
port 15 nsew ground bidirectional
rlabel metal2 s 2410 0 2466 800 6 xi0[0]
port 16 nsew signal input
rlabel metal2 s 9034 0 9090 800 6 xi0[1]
port 17 nsew signal input
rlabel metal2 s 15658 0 15714 800 6 xi0[2]
port 18 nsew signal input
rlabel metal2 s 22282 0 22338 800 6 xi0[3]
port 19 nsew signal input
rlabel metal2 s 4066 0 4122 800 6 xi1[0]
port 20 nsew signal input
rlabel metal2 s 10690 0 10746 800 6 xi1[1]
port 21 nsew signal input
rlabel metal2 s 17314 0 17370 800 6 xi1[2]
port 22 nsew signal input
rlabel metal2 s 23938 0 23994 800 6 xi1[3]
port 23 nsew signal input
rlabel metal2 s 5722 0 5778 800 6 xi2[0]
port 24 nsew signal input
rlabel metal2 s 12346 0 12402 800 6 xi2[1]
port 25 nsew signal input
rlabel metal2 s 18970 0 19026 800 6 xi2[2]
port 26 nsew signal input
rlabel metal2 s 25594 0 25650 800 6 xi2[3]
port 27 nsew signal input
rlabel metal2 s 7378 0 7434 800 6 xi3[0]
port 28 nsew signal input
rlabel metal2 s 14002 0 14058 800 6 xi3[1]
port 29 nsew signal input
rlabel metal2 s 20626 0 20682 800 6 xi3[2]
port 30 nsew signal input
rlabel metal2 s 27250 0 27306 800 6 xi3[3]
port 31 nsew signal input
rlabel metal2 s 1582 0 1638 800 6 xr0[0]
port 32 nsew signal input
rlabel metal2 s 8206 0 8262 800 6 xr0[1]
port 33 nsew signal input
rlabel metal2 s 14830 0 14886 800 6 xr0[2]
port 34 nsew signal input
rlabel metal2 s 21454 0 21510 800 6 xr0[3]
port 35 nsew signal input
rlabel metal2 s 3238 0 3294 800 6 xr1[0]
port 36 nsew signal input
rlabel metal2 s 9862 0 9918 800 6 xr1[1]
port 37 nsew signal input
rlabel metal2 s 16486 0 16542 800 6 xr1[2]
port 38 nsew signal input
rlabel metal2 s 23110 0 23166 800 6 xr1[3]
port 39 nsew signal input
rlabel metal2 s 4894 0 4950 800 6 xr2[0]
port 40 nsew signal input
rlabel metal2 s 11518 0 11574 800 6 xr2[1]
port 41 nsew signal input
rlabel metal2 s 18142 0 18198 800 6 xr2[2]
port 42 nsew signal input
rlabel metal2 s 24766 0 24822 800 6 xr2[3]
port 43 nsew signal input
rlabel metal2 s 6550 0 6606 800 6 xr3[0]
port 44 nsew signal input
rlabel metal2 s 13174 0 13230 800 6 xr3[1]
port 45 nsew signal input
rlabel metal2 s 19798 0 19854 800 6 xr3[2]
port 46 nsew signal input
rlabel metal2 s 26422 0 26478 800 6 xr3[3]
port 47 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 36400 38800
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 500560
string GDS_FILE /home/guanyanlye/unic-cass/caravel_tutorial/UNICCASS_copy/openlane/R4_butter/runs/23_11_09_00_02/results/signoff/R4_butter.magic.gds
string GDS_START 80640
<< end >>

