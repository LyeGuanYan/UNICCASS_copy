VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO R4_butter
  CLASS BLOCK ;
  FOREIGN R4_butter ;
  ORIGIN 0.000 0.000 ;
  SIZE 182.000 BY 194.000 ;
  PIN Xio[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 178.000 46.280 182.000 46.880 ;
    END
  END Xio[0]
  PIN Xio[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 178.000 93.880 182.000 94.480 ;
    END
  END Xio[1]
  PIN Xio[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 178.000 141.480 182.000 142.080 ;
    END
  END Xio[2]
  PIN Xio[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 178.000 189.080 182.000 189.680 ;
    END
  END Xio[3]
  PIN Xro[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 178.000 41.520 182.000 42.120 ;
    END
  END Xro[0]
  PIN Xro[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 178.000 89.120 182.000 89.720 ;
    END
  END Xro[1]
  PIN Xro[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 178.000 136.720 182.000 137.320 ;
    END
  END Xro[2]
  PIN Xro[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 178.000 184.320 182.000 184.920 ;
    END
  END Xro[3]
  PIN c1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 161.200 4.000 161.800 ;
    END
  END c1
  PIN c2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 96.600 4.000 97.200 ;
    END
  END c2
  PIN c3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 32.000 4.000 32.600 ;
    END
  END c3
  PIN la_oenb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 12.050 0.000 12.330 4.000 ;
    END
  END la_oenb[0]
  PIN la_oenb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 34.590 0.000 34.870 4.000 ;
    END
  END la_oenb[1]
  PIN la_oenb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 57.130 0.000 57.410 4.000 ;
    END
  END la_oenb[2]
  PIN la_oenb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 79.670 0.000 79.950 4.000 ;
    END
  END la_oenb[3]
  PIN la_oenb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 102.210 0.000 102.490 4.000 ;
    END
  END la_oenb[4]
  PIN la_oenb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 124.750 0.000 125.030 4.000 ;
    END
  END la_oenb[5]
  PIN la_oenb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 147.290 0.000 147.570 4.000 ;
    END
  END la_oenb[6]
  PIN la_oenb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 169.830 0.000 170.110 4.000 ;
    END
  END la_oenb[7]
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 182.480 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 182.480 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 182.480 ;
    END
  END vssd1
  PIN xi0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 178.000 8.200 182.000 8.800 ;
    END
  END xi0[0]
  PIN xi0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 178.000 55.800 182.000 56.400 ;
    END
  END xi0[1]
  PIN xi0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 178.000 103.400 182.000 104.000 ;
    END
  END xi0[2]
  PIN xi0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 178.000 151.000 182.000 151.600 ;
    END
  END xi0[3]
  PIN xi1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 178.000 17.720 182.000 18.320 ;
    END
  END xi1[0]
  PIN xi1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 178.000 65.320 182.000 65.920 ;
    END
  END xi1[1]
  PIN xi1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 178.000 112.920 182.000 113.520 ;
    END
  END xi1[2]
  PIN xi1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 178.000 160.520 182.000 161.120 ;
    END
  END xi1[3]
  PIN xi2[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 178.000 27.240 182.000 27.840 ;
    END
  END xi2[0]
  PIN xi2[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 178.000 74.840 182.000 75.440 ;
    END
  END xi2[1]
  PIN xi2[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 178.000 122.440 182.000 123.040 ;
    END
  END xi2[2]
  PIN xi2[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 178.000 170.040 182.000 170.640 ;
    END
  END xi2[3]
  PIN xi3[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 178.000 36.760 182.000 37.360 ;
    END
  END xi3[0]
  PIN xi3[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 178.000 84.360 182.000 84.960 ;
    END
  END xi3[1]
  PIN xi3[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 178.000 131.960 182.000 132.560 ;
    END
  END xi3[2]
  PIN xi3[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 178.000 179.560 182.000 180.160 ;
    END
  END xi3[3]
  PIN xr0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 178.000 3.440 182.000 4.040 ;
    END
  END xr0[0]
  PIN xr0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 178.000 51.040 182.000 51.640 ;
    END
  END xr0[1]
  PIN xr0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 178.000 98.640 182.000 99.240 ;
    END
  END xr0[2]
  PIN xr0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 178.000 146.240 182.000 146.840 ;
    END
  END xr0[3]
  PIN xr1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 178.000 12.960 182.000 13.560 ;
    END
  END xr1[0]
  PIN xr1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 178.000 60.560 182.000 61.160 ;
    END
  END xr1[1]
  PIN xr1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 178.000 108.160 182.000 108.760 ;
    END
  END xr1[2]
  PIN xr1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 178.000 155.760 182.000 156.360 ;
    END
  END xr1[3]
  PIN xr2[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 178.000 22.480 182.000 23.080 ;
    END
  END xr2[0]
  PIN xr2[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 178.000 70.080 182.000 70.680 ;
    END
  END xr2[1]
  PIN xr2[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 178.000 117.680 182.000 118.280 ;
    END
  END xr2[2]
  PIN xr2[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 178.000 165.280 182.000 165.880 ;
    END
  END xr2[3]
  PIN xr3[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 178.000 32.000 182.000 32.600 ;
    END
  END xr3[0]
  PIN xr3[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 178.000 79.600 182.000 80.200 ;
    END
  END xr3[1]
  PIN xr3[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 178.000 127.200 182.000 127.800 ;
    END
  END xr3[2]
  PIN xr3[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 178.000 174.800 182.000 175.400 ;
    END
  END xr3[3]
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 176.180 182.325 ;
      LAYER met1 ;
        RECT 4.670 10.640 177.490 182.480 ;
      LAYER met2 ;
        RECT 4.690 4.280 177.470 189.565 ;
        RECT 4.690 3.555 11.770 4.280 ;
        RECT 12.610 3.555 34.310 4.280 ;
        RECT 35.150 3.555 56.850 4.280 ;
        RECT 57.690 3.555 79.390 4.280 ;
        RECT 80.230 3.555 101.930 4.280 ;
        RECT 102.770 3.555 124.470 4.280 ;
        RECT 125.310 3.555 147.010 4.280 ;
        RECT 147.850 3.555 169.550 4.280 ;
        RECT 170.390 3.555 177.470 4.280 ;
      LAYER met3 ;
        RECT 4.000 188.680 177.600 189.545 ;
        RECT 4.000 185.320 178.000 188.680 ;
        RECT 4.000 183.920 177.600 185.320 ;
        RECT 4.000 180.560 178.000 183.920 ;
        RECT 4.000 179.160 177.600 180.560 ;
        RECT 4.000 175.800 178.000 179.160 ;
        RECT 4.000 174.400 177.600 175.800 ;
        RECT 4.000 171.040 178.000 174.400 ;
        RECT 4.000 169.640 177.600 171.040 ;
        RECT 4.000 166.280 178.000 169.640 ;
        RECT 4.000 164.880 177.600 166.280 ;
        RECT 4.000 162.200 178.000 164.880 ;
        RECT 4.400 161.520 178.000 162.200 ;
        RECT 4.400 160.800 177.600 161.520 ;
        RECT 4.000 160.120 177.600 160.800 ;
        RECT 4.000 156.760 178.000 160.120 ;
        RECT 4.000 155.360 177.600 156.760 ;
        RECT 4.000 152.000 178.000 155.360 ;
        RECT 4.000 150.600 177.600 152.000 ;
        RECT 4.000 147.240 178.000 150.600 ;
        RECT 4.000 145.840 177.600 147.240 ;
        RECT 4.000 142.480 178.000 145.840 ;
        RECT 4.000 141.080 177.600 142.480 ;
        RECT 4.000 137.720 178.000 141.080 ;
        RECT 4.000 136.320 177.600 137.720 ;
        RECT 4.000 132.960 178.000 136.320 ;
        RECT 4.000 131.560 177.600 132.960 ;
        RECT 4.000 128.200 178.000 131.560 ;
        RECT 4.000 126.800 177.600 128.200 ;
        RECT 4.000 123.440 178.000 126.800 ;
        RECT 4.000 122.040 177.600 123.440 ;
        RECT 4.000 118.680 178.000 122.040 ;
        RECT 4.000 117.280 177.600 118.680 ;
        RECT 4.000 113.920 178.000 117.280 ;
        RECT 4.000 112.520 177.600 113.920 ;
        RECT 4.000 109.160 178.000 112.520 ;
        RECT 4.000 107.760 177.600 109.160 ;
        RECT 4.000 104.400 178.000 107.760 ;
        RECT 4.000 103.000 177.600 104.400 ;
        RECT 4.000 99.640 178.000 103.000 ;
        RECT 4.000 98.240 177.600 99.640 ;
        RECT 4.000 97.600 178.000 98.240 ;
        RECT 4.400 96.200 178.000 97.600 ;
        RECT 4.000 94.880 178.000 96.200 ;
        RECT 4.000 93.480 177.600 94.880 ;
        RECT 4.000 90.120 178.000 93.480 ;
        RECT 4.000 88.720 177.600 90.120 ;
        RECT 4.000 85.360 178.000 88.720 ;
        RECT 4.000 83.960 177.600 85.360 ;
        RECT 4.000 80.600 178.000 83.960 ;
        RECT 4.000 79.200 177.600 80.600 ;
        RECT 4.000 75.840 178.000 79.200 ;
        RECT 4.000 74.440 177.600 75.840 ;
        RECT 4.000 71.080 178.000 74.440 ;
        RECT 4.000 69.680 177.600 71.080 ;
        RECT 4.000 66.320 178.000 69.680 ;
        RECT 4.000 64.920 177.600 66.320 ;
        RECT 4.000 61.560 178.000 64.920 ;
        RECT 4.000 60.160 177.600 61.560 ;
        RECT 4.000 56.800 178.000 60.160 ;
        RECT 4.000 55.400 177.600 56.800 ;
        RECT 4.000 52.040 178.000 55.400 ;
        RECT 4.000 50.640 177.600 52.040 ;
        RECT 4.000 47.280 178.000 50.640 ;
        RECT 4.000 45.880 177.600 47.280 ;
        RECT 4.000 42.520 178.000 45.880 ;
        RECT 4.000 41.120 177.600 42.520 ;
        RECT 4.000 37.760 178.000 41.120 ;
        RECT 4.000 36.360 177.600 37.760 ;
        RECT 4.000 33.000 178.000 36.360 ;
        RECT 4.400 31.600 177.600 33.000 ;
        RECT 4.000 28.240 178.000 31.600 ;
        RECT 4.000 26.840 177.600 28.240 ;
        RECT 4.000 23.480 178.000 26.840 ;
        RECT 4.000 22.080 177.600 23.480 ;
        RECT 4.000 18.720 178.000 22.080 ;
        RECT 4.000 17.320 177.600 18.720 ;
        RECT 4.000 13.960 178.000 17.320 ;
        RECT 4.000 12.560 177.600 13.960 ;
        RECT 4.000 9.200 178.000 12.560 ;
        RECT 4.000 7.800 177.600 9.200 ;
        RECT 4.000 4.440 178.000 7.800 ;
        RECT 4.000 3.575 177.600 4.440 ;
  END
END R4_butter
END LIBRARY

