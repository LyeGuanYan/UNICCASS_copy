magic
tech sky130A
magscale 1 2
timestamp 1696211632
<< obsli1 >>
rect 1104 2159 558808 349809
<< obsm1 >>
rect 934 2128 558808 349840
<< obsm2 >>
rect 938 2139 558422 349829
<< metal3 >>
rect 559200 345584 560000 345704
rect 559200 336880 560000 337000
rect 559200 328176 560000 328296
rect 559200 319472 560000 319592
rect 559200 310768 560000 310888
rect 559200 302064 560000 302184
rect 559200 293360 560000 293480
rect 0 293088 800 293208
rect 559200 284656 560000 284776
rect 559200 275952 560000 276072
rect 559200 267248 560000 267368
rect 559200 258544 560000 258664
rect 559200 249840 560000 249960
rect 559200 241136 560000 241256
rect 559200 232432 560000 232552
rect 559200 223728 560000 223848
rect 559200 215024 560000 215144
rect 559200 206320 560000 206440
rect 559200 197616 560000 197736
rect 559200 188912 560000 189032
rect 559200 180208 560000 180328
rect 0 175856 800 175976
rect 559200 171504 560000 171624
rect 559200 162800 560000 162920
rect 559200 154096 560000 154216
rect 559200 145392 560000 145512
rect 559200 136688 560000 136808
rect 559200 127984 560000 128104
rect 559200 119280 560000 119400
rect 559200 110576 560000 110696
rect 559200 101872 560000 101992
rect 559200 93168 560000 93288
rect 559200 84464 560000 84584
rect 559200 75760 560000 75880
rect 559200 67056 560000 67176
rect 0 58624 800 58744
rect 559200 58352 560000 58472
rect 559200 49648 560000 49768
rect 559200 40944 560000 41064
rect 559200 32240 560000 32360
rect 559200 23536 560000 23656
rect 559200 14832 560000 14952
rect 559200 6128 560000 6248
<< obsm3 >>
rect 800 345784 559200 349825
rect 800 345504 559120 345784
rect 800 337080 559200 345504
rect 800 336800 559120 337080
rect 800 328376 559200 336800
rect 800 328096 559120 328376
rect 800 319672 559200 328096
rect 800 319392 559120 319672
rect 800 310968 559200 319392
rect 800 310688 559120 310968
rect 800 302264 559200 310688
rect 800 301984 559120 302264
rect 800 293560 559200 301984
rect 800 293288 559120 293560
rect 880 293280 559120 293288
rect 880 293008 559200 293280
rect 800 284856 559200 293008
rect 800 284576 559120 284856
rect 800 276152 559200 284576
rect 800 275872 559120 276152
rect 800 267448 559200 275872
rect 800 267168 559120 267448
rect 800 258744 559200 267168
rect 800 258464 559120 258744
rect 800 250040 559200 258464
rect 800 249760 559120 250040
rect 800 241336 559200 249760
rect 800 241056 559120 241336
rect 800 232632 559200 241056
rect 800 232352 559120 232632
rect 800 223928 559200 232352
rect 800 223648 559120 223928
rect 800 215224 559200 223648
rect 800 214944 559120 215224
rect 800 206520 559200 214944
rect 800 206240 559120 206520
rect 800 197816 559200 206240
rect 800 197536 559120 197816
rect 800 189112 559200 197536
rect 800 188832 559120 189112
rect 800 180408 559200 188832
rect 800 180128 559120 180408
rect 800 176056 559200 180128
rect 880 175776 559200 176056
rect 800 171704 559200 175776
rect 800 171424 559120 171704
rect 800 163000 559200 171424
rect 800 162720 559120 163000
rect 800 154296 559200 162720
rect 800 154016 559120 154296
rect 800 145592 559200 154016
rect 800 145312 559120 145592
rect 800 136888 559200 145312
rect 800 136608 559120 136888
rect 800 128184 559200 136608
rect 800 127904 559120 128184
rect 800 119480 559200 127904
rect 800 119200 559120 119480
rect 800 110776 559200 119200
rect 800 110496 559120 110776
rect 800 102072 559200 110496
rect 800 101792 559120 102072
rect 800 93368 559200 101792
rect 800 93088 559120 93368
rect 800 84664 559200 93088
rect 800 84384 559120 84664
rect 800 75960 559200 84384
rect 800 75680 559120 75960
rect 800 67256 559200 75680
rect 800 66976 559120 67256
rect 800 58824 559200 66976
rect 880 58552 559200 58824
rect 880 58544 559120 58552
rect 800 58272 559120 58544
rect 800 49848 559200 58272
rect 800 49568 559120 49848
rect 800 41144 559200 49568
rect 800 40864 559120 41144
rect 800 32440 559200 40864
rect 800 32160 559120 32440
rect 800 23736 559200 32160
rect 800 23456 559120 23736
rect 800 15032 559200 23456
rect 800 14752 559120 15032
rect 800 6328 559200 14752
rect 800 6048 559120 6328
rect 800 2143 559200 6048
<< metal4 >>
rect 4208 2128 4528 349840
rect 19568 2128 19888 349840
rect 34928 2128 35248 349840
rect 50288 2128 50608 349840
rect 65648 2128 65968 349840
rect 81008 2128 81328 349840
rect 96368 2128 96688 349840
rect 111728 2128 112048 349840
rect 127088 2128 127408 349840
rect 142448 2128 142768 349840
rect 157808 2128 158128 349840
rect 173168 2128 173488 349840
rect 188528 2128 188848 349840
rect 203888 2128 204208 349840
rect 219248 2128 219568 349840
rect 234608 2128 234928 349840
rect 249968 2128 250288 349840
rect 265328 2128 265648 349840
rect 280688 2128 281008 349840
rect 296048 2128 296368 349840
rect 311408 2128 311728 349840
rect 326768 2128 327088 349840
rect 342128 2128 342448 349840
rect 357488 2128 357808 349840
rect 372848 2128 373168 349840
rect 388208 2128 388528 349840
rect 403568 2128 403888 349840
rect 418928 2128 419248 349840
rect 434288 2128 434608 349840
rect 449648 2128 449968 349840
rect 465008 2128 465328 349840
rect 480368 2128 480688 349840
rect 495728 2128 496048 349840
rect 511088 2128 511408 349840
rect 526448 2128 526768 349840
rect 541808 2128 542128 349840
rect 557168 2128 557488 349840
<< labels >>
rlabel metal3 s 559200 84464 560000 84584 6 Xio[0]
port 1 nsew signal output
rlabel metal3 s 559200 171504 560000 171624 6 Xio[1]
port 2 nsew signal output
rlabel metal3 s 559200 258544 560000 258664 6 Xio[2]
port 3 nsew signal output
rlabel metal3 s 559200 345584 560000 345704 6 Xio[3]
port 4 nsew signal output
rlabel metal3 s 559200 75760 560000 75880 6 Xro[0]
port 5 nsew signal output
rlabel metal3 s 559200 162800 560000 162920 6 Xro[1]
port 6 nsew signal output
rlabel metal3 s 559200 249840 560000 249960 6 Xro[2]
port 7 nsew signal output
rlabel metal3 s 559200 336880 560000 337000 6 Xro[3]
port 8 nsew signal output
rlabel metal3 s 0 293088 800 293208 6 c1
port 9 nsew signal input
rlabel metal3 s 0 175856 800 175976 6 c2
port 10 nsew signal input
rlabel metal3 s 0 58624 800 58744 6 c3
port 11 nsew signal input
rlabel metal4 s 4208 2128 4528 349840 6 vccd1
port 12 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 349840 6 vccd1
port 12 nsew power bidirectional
rlabel metal4 s 65648 2128 65968 349840 6 vccd1
port 12 nsew power bidirectional
rlabel metal4 s 96368 2128 96688 349840 6 vccd1
port 12 nsew power bidirectional
rlabel metal4 s 127088 2128 127408 349840 6 vccd1
port 12 nsew power bidirectional
rlabel metal4 s 157808 2128 158128 349840 6 vccd1
port 12 nsew power bidirectional
rlabel metal4 s 188528 2128 188848 349840 6 vccd1
port 12 nsew power bidirectional
rlabel metal4 s 219248 2128 219568 349840 6 vccd1
port 12 nsew power bidirectional
rlabel metal4 s 249968 2128 250288 349840 6 vccd1
port 12 nsew power bidirectional
rlabel metal4 s 280688 2128 281008 349840 6 vccd1
port 12 nsew power bidirectional
rlabel metal4 s 311408 2128 311728 349840 6 vccd1
port 12 nsew power bidirectional
rlabel metal4 s 342128 2128 342448 349840 6 vccd1
port 12 nsew power bidirectional
rlabel metal4 s 372848 2128 373168 349840 6 vccd1
port 12 nsew power bidirectional
rlabel metal4 s 403568 2128 403888 349840 6 vccd1
port 12 nsew power bidirectional
rlabel metal4 s 434288 2128 434608 349840 6 vccd1
port 12 nsew power bidirectional
rlabel metal4 s 465008 2128 465328 349840 6 vccd1
port 12 nsew power bidirectional
rlabel metal4 s 495728 2128 496048 349840 6 vccd1
port 12 nsew power bidirectional
rlabel metal4 s 526448 2128 526768 349840 6 vccd1
port 12 nsew power bidirectional
rlabel metal4 s 557168 2128 557488 349840 6 vccd1
port 12 nsew power bidirectional
rlabel metal4 s 19568 2128 19888 349840 6 vssd1
port 13 nsew ground bidirectional
rlabel metal4 s 50288 2128 50608 349840 6 vssd1
port 13 nsew ground bidirectional
rlabel metal4 s 81008 2128 81328 349840 6 vssd1
port 13 nsew ground bidirectional
rlabel metal4 s 111728 2128 112048 349840 6 vssd1
port 13 nsew ground bidirectional
rlabel metal4 s 142448 2128 142768 349840 6 vssd1
port 13 nsew ground bidirectional
rlabel metal4 s 173168 2128 173488 349840 6 vssd1
port 13 nsew ground bidirectional
rlabel metal4 s 203888 2128 204208 349840 6 vssd1
port 13 nsew ground bidirectional
rlabel metal4 s 234608 2128 234928 349840 6 vssd1
port 13 nsew ground bidirectional
rlabel metal4 s 265328 2128 265648 349840 6 vssd1
port 13 nsew ground bidirectional
rlabel metal4 s 296048 2128 296368 349840 6 vssd1
port 13 nsew ground bidirectional
rlabel metal4 s 326768 2128 327088 349840 6 vssd1
port 13 nsew ground bidirectional
rlabel metal4 s 357488 2128 357808 349840 6 vssd1
port 13 nsew ground bidirectional
rlabel metal4 s 388208 2128 388528 349840 6 vssd1
port 13 nsew ground bidirectional
rlabel metal4 s 418928 2128 419248 349840 6 vssd1
port 13 nsew ground bidirectional
rlabel metal4 s 449648 2128 449968 349840 6 vssd1
port 13 nsew ground bidirectional
rlabel metal4 s 480368 2128 480688 349840 6 vssd1
port 13 nsew ground bidirectional
rlabel metal4 s 511088 2128 511408 349840 6 vssd1
port 13 nsew ground bidirectional
rlabel metal4 s 541808 2128 542128 349840 6 vssd1
port 13 nsew ground bidirectional
rlabel metal3 s 559200 14832 560000 14952 6 xi0[0]
port 14 nsew signal input
rlabel metal3 s 559200 101872 560000 101992 6 xi0[1]
port 15 nsew signal input
rlabel metal3 s 559200 188912 560000 189032 6 xi0[2]
port 16 nsew signal input
rlabel metal3 s 559200 275952 560000 276072 6 xi0[3]
port 17 nsew signal input
rlabel metal3 s 559200 32240 560000 32360 6 xi1[0]
port 18 nsew signal input
rlabel metal3 s 559200 119280 560000 119400 6 xi1[1]
port 19 nsew signal input
rlabel metal3 s 559200 206320 560000 206440 6 xi1[2]
port 20 nsew signal input
rlabel metal3 s 559200 293360 560000 293480 6 xi1[3]
port 21 nsew signal input
rlabel metal3 s 559200 49648 560000 49768 6 xi2[0]
port 22 nsew signal input
rlabel metal3 s 559200 136688 560000 136808 6 xi2[1]
port 23 nsew signal input
rlabel metal3 s 559200 223728 560000 223848 6 xi2[2]
port 24 nsew signal input
rlabel metal3 s 559200 310768 560000 310888 6 xi2[3]
port 25 nsew signal input
rlabel metal3 s 559200 67056 560000 67176 6 xi3[0]
port 26 nsew signal input
rlabel metal3 s 559200 154096 560000 154216 6 xi3[1]
port 27 nsew signal input
rlabel metal3 s 559200 241136 560000 241256 6 xi3[2]
port 28 nsew signal input
rlabel metal3 s 559200 328176 560000 328296 6 xi3[3]
port 29 nsew signal input
rlabel metal3 s 559200 6128 560000 6248 6 xr0[0]
port 30 nsew signal input
rlabel metal3 s 559200 93168 560000 93288 6 xr0[1]
port 31 nsew signal input
rlabel metal3 s 559200 180208 560000 180328 6 xr0[2]
port 32 nsew signal input
rlabel metal3 s 559200 267248 560000 267368 6 xr0[3]
port 33 nsew signal input
rlabel metal3 s 559200 23536 560000 23656 6 xr1[0]
port 34 nsew signal input
rlabel metal3 s 559200 110576 560000 110696 6 xr1[1]
port 35 nsew signal input
rlabel metal3 s 559200 197616 560000 197736 6 xr1[2]
port 36 nsew signal input
rlabel metal3 s 559200 284656 560000 284776 6 xr1[3]
port 37 nsew signal input
rlabel metal3 s 559200 40944 560000 41064 6 xr2[0]
port 38 nsew signal input
rlabel metal3 s 559200 127984 560000 128104 6 xr2[1]
port 39 nsew signal input
rlabel metal3 s 559200 215024 560000 215144 6 xr2[2]
port 40 nsew signal input
rlabel metal3 s 559200 302064 560000 302184 6 xr2[3]
port 41 nsew signal input
rlabel metal3 s 559200 58352 560000 58472 6 xr3[0]
port 42 nsew signal input
rlabel metal3 s 559200 145392 560000 145512 6 xr3[1]
port 43 nsew signal input
rlabel metal3 s 559200 232432 560000 232552 6 xr3[2]
port 44 nsew signal input
rlabel metal3 s 559200 319472 560000 319592 6 xr3[3]
port 45 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 560000 352000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 50688130
string GDS_FILE /home/guanyanlye/unic-cass/caravel_tutorial/caravel_uniccas_example/openlane/R4_butter/runs/23_10_02_09_44/results/signoff/R4_butter.magic.gds
string GDS_START 96716
<< end >>

