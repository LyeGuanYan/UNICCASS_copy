VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO R4_butter
  CLASS BLOCK ;
  FOREIGN R4_butter ;
  ORIGIN 0.000 0.000 ;
  SIZE 2800.000 BY 1760.000 ;
  PIN Xio[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2796.000 422.320 2800.000 422.920 ;
    END
  END Xio[0]
  PIN Xio[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2796.000 857.520 2800.000 858.120 ;
    END
  END Xio[1]
  PIN Xio[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2796.000 1292.720 2800.000 1293.320 ;
    END
  END Xio[2]
  PIN Xio[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2796.000 1727.920 2800.000 1728.520 ;
    END
  END Xio[3]
  PIN Xro[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2796.000 378.800 2800.000 379.400 ;
    END
  END Xro[0]
  PIN Xro[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2796.000 814.000 2800.000 814.600 ;
    END
  END Xro[1]
  PIN Xro[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2796.000 1249.200 2800.000 1249.800 ;
    END
  END Xro[2]
  PIN Xro[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2796.000 1684.400 2800.000 1685.000 ;
    END
  END Xro[3]
  PIN c1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1465.440 4.000 1466.040 ;
    END
  END c1
  PIN c2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 879.280 4.000 879.880 ;
    END
  END c2
  PIN c3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 293.120 4.000 293.720 ;
    END
  END c3
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 481.840 10.640 483.440 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 635.440 10.640 637.040 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 789.040 10.640 790.640 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 942.640 10.640 944.240 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 1096.240 10.640 1097.840 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 1249.840 10.640 1251.440 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 1403.440 10.640 1405.040 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 1557.040 10.640 1558.640 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 1710.640 10.640 1712.240 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 1864.240 10.640 1865.840 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 2017.840 10.640 2019.440 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 2171.440 10.640 2173.040 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 2325.040 10.640 2326.640 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 2478.640 10.640 2480.240 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 2632.240 10.640 2633.840 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 2785.840 10.640 2787.440 1749.200 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 405.040 10.640 406.640 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 558.640 10.640 560.240 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 712.240 10.640 713.840 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 865.840 10.640 867.440 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 1019.440 10.640 1021.040 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 1173.040 10.640 1174.640 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 1326.640 10.640 1328.240 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 1480.240 10.640 1481.840 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 1633.840 10.640 1635.440 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 1787.440 10.640 1789.040 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 1941.040 10.640 1942.640 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 2094.640 10.640 2096.240 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 2248.240 10.640 2249.840 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 2401.840 10.640 2403.440 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 2555.440 10.640 2557.040 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 2709.040 10.640 2710.640 1749.200 ;
    END
  END vssd1
  PIN xi0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2796.000 74.160 2800.000 74.760 ;
    END
  END xi0[0]
  PIN xi0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2796.000 509.360 2800.000 509.960 ;
    END
  END xi0[1]
  PIN xi0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2796.000 944.560 2800.000 945.160 ;
    END
  END xi0[2]
  PIN xi0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2796.000 1379.760 2800.000 1380.360 ;
    END
  END xi0[3]
  PIN xi1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2796.000 161.200 2800.000 161.800 ;
    END
  END xi1[0]
  PIN xi1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2796.000 596.400 2800.000 597.000 ;
    END
  END xi1[1]
  PIN xi1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2796.000 1031.600 2800.000 1032.200 ;
    END
  END xi1[2]
  PIN xi1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2796.000 1466.800 2800.000 1467.400 ;
    END
  END xi1[3]
  PIN xi2[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2796.000 248.240 2800.000 248.840 ;
    END
  END xi2[0]
  PIN xi2[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2796.000 683.440 2800.000 684.040 ;
    END
  END xi2[1]
  PIN xi2[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2796.000 1118.640 2800.000 1119.240 ;
    END
  END xi2[2]
  PIN xi2[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2796.000 1553.840 2800.000 1554.440 ;
    END
  END xi2[3]
  PIN xi3[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2796.000 335.280 2800.000 335.880 ;
    END
  END xi3[0]
  PIN xi3[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2796.000 770.480 2800.000 771.080 ;
    END
  END xi3[1]
  PIN xi3[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2796.000 1205.680 2800.000 1206.280 ;
    END
  END xi3[2]
  PIN xi3[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2796.000 1640.880 2800.000 1641.480 ;
    END
  END xi3[3]
  PIN xr0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2796.000 30.640 2800.000 31.240 ;
    END
  END xr0[0]
  PIN xr0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2796.000 465.840 2800.000 466.440 ;
    END
  END xr0[1]
  PIN xr0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2796.000 901.040 2800.000 901.640 ;
    END
  END xr0[2]
  PIN xr0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2796.000 1336.240 2800.000 1336.840 ;
    END
  END xr0[3]
  PIN xr1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2796.000 117.680 2800.000 118.280 ;
    END
  END xr1[0]
  PIN xr1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2796.000 552.880 2800.000 553.480 ;
    END
  END xr1[1]
  PIN xr1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2796.000 988.080 2800.000 988.680 ;
    END
  END xr1[2]
  PIN xr1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2796.000 1423.280 2800.000 1423.880 ;
    END
  END xr1[3]
  PIN xr2[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2796.000 204.720 2800.000 205.320 ;
    END
  END xr2[0]
  PIN xr2[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2796.000 639.920 2800.000 640.520 ;
    END
  END xr2[1]
  PIN xr2[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2796.000 1075.120 2800.000 1075.720 ;
    END
  END xr2[2]
  PIN xr2[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2796.000 1510.320 2800.000 1510.920 ;
    END
  END xr2[3]
  PIN xr3[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2796.000 291.760 2800.000 292.360 ;
    END
  END xr3[0]
  PIN xr3[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2796.000 726.960 2800.000 727.560 ;
    END
  END xr3[1]
  PIN xr3[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2796.000 1162.160 2800.000 1162.760 ;
    END
  END xr3[2]
  PIN xr3[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2796.000 1597.360 2800.000 1597.960 ;
    END
  END xr3[3]
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 2794.040 1749.045 ;
      LAYER met1 ;
        RECT 4.670 10.640 2794.040 1749.200 ;
      LAYER met2 ;
        RECT 4.690 10.695 2792.110 1749.145 ;
      LAYER met3 ;
        RECT 4.000 1728.920 2796.000 1749.125 ;
        RECT 4.000 1727.520 2795.600 1728.920 ;
        RECT 4.000 1685.400 2796.000 1727.520 ;
        RECT 4.000 1684.000 2795.600 1685.400 ;
        RECT 4.000 1641.880 2796.000 1684.000 ;
        RECT 4.000 1640.480 2795.600 1641.880 ;
        RECT 4.000 1598.360 2796.000 1640.480 ;
        RECT 4.000 1596.960 2795.600 1598.360 ;
        RECT 4.000 1554.840 2796.000 1596.960 ;
        RECT 4.000 1553.440 2795.600 1554.840 ;
        RECT 4.000 1511.320 2796.000 1553.440 ;
        RECT 4.000 1509.920 2795.600 1511.320 ;
        RECT 4.000 1467.800 2796.000 1509.920 ;
        RECT 4.000 1466.440 2795.600 1467.800 ;
        RECT 4.400 1466.400 2795.600 1466.440 ;
        RECT 4.400 1465.040 2796.000 1466.400 ;
        RECT 4.000 1424.280 2796.000 1465.040 ;
        RECT 4.000 1422.880 2795.600 1424.280 ;
        RECT 4.000 1380.760 2796.000 1422.880 ;
        RECT 4.000 1379.360 2795.600 1380.760 ;
        RECT 4.000 1337.240 2796.000 1379.360 ;
        RECT 4.000 1335.840 2795.600 1337.240 ;
        RECT 4.000 1293.720 2796.000 1335.840 ;
        RECT 4.000 1292.320 2795.600 1293.720 ;
        RECT 4.000 1250.200 2796.000 1292.320 ;
        RECT 4.000 1248.800 2795.600 1250.200 ;
        RECT 4.000 1206.680 2796.000 1248.800 ;
        RECT 4.000 1205.280 2795.600 1206.680 ;
        RECT 4.000 1163.160 2796.000 1205.280 ;
        RECT 4.000 1161.760 2795.600 1163.160 ;
        RECT 4.000 1119.640 2796.000 1161.760 ;
        RECT 4.000 1118.240 2795.600 1119.640 ;
        RECT 4.000 1076.120 2796.000 1118.240 ;
        RECT 4.000 1074.720 2795.600 1076.120 ;
        RECT 4.000 1032.600 2796.000 1074.720 ;
        RECT 4.000 1031.200 2795.600 1032.600 ;
        RECT 4.000 989.080 2796.000 1031.200 ;
        RECT 4.000 987.680 2795.600 989.080 ;
        RECT 4.000 945.560 2796.000 987.680 ;
        RECT 4.000 944.160 2795.600 945.560 ;
        RECT 4.000 902.040 2796.000 944.160 ;
        RECT 4.000 900.640 2795.600 902.040 ;
        RECT 4.000 880.280 2796.000 900.640 ;
        RECT 4.400 878.880 2796.000 880.280 ;
        RECT 4.000 858.520 2796.000 878.880 ;
        RECT 4.000 857.120 2795.600 858.520 ;
        RECT 4.000 815.000 2796.000 857.120 ;
        RECT 4.000 813.600 2795.600 815.000 ;
        RECT 4.000 771.480 2796.000 813.600 ;
        RECT 4.000 770.080 2795.600 771.480 ;
        RECT 4.000 727.960 2796.000 770.080 ;
        RECT 4.000 726.560 2795.600 727.960 ;
        RECT 4.000 684.440 2796.000 726.560 ;
        RECT 4.000 683.040 2795.600 684.440 ;
        RECT 4.000 640.920 2796.000 683.040 ;
        RECT 4.000 639.520 2795.600 640.920 ;
        RECT 4.000 597.400 2796.000 639.520 ;
        RECT 4.000 596.000 2795.600 597.400 ;
        RECT 4.000 553.880 2796.000 596.000 ;
        RECT 4.000 552.480 2795.600 553.880 ;
        RECT 4.000 510.360 2796.000 552.480 ;
        RECT 4.000 508.960 2795.600 510.360 ;
        RECT 4.000 466.840 2796.000 508.960 ;
        RECT 4.000 465.440 2795.600 466.840 ;
        RECT 4.000 423.320 2796.000 465.440 ;
        RECT 4.000 421.920 2795.600 423.320 ;
        RECT 4.000 379.800 2796.000 421.920 ;
        RECT 4.000 378.400 2795.600 379.800 ;
        RECT 4.000 336.280 2796.000 378.400 ;
        RECT 4.000 334.880 2795.600 336.280 ;
        RECT 4.000 294.120 2796.000 334.880 ;
        RECT 4.400 292.760 2796.000 294.120 ;
        RECT 4.400 292.720 2795.600 292.760 ;
        RECT 4.000 291.360 2795.600 292.720 ;
        RECT 4.000 249.240 2796.000 291.360 ;
        RECT 4.000 247.840 2795.600 249.240 ;
        RECT 4.000 205.720 2796.000 247.840 ;
        RECT 4.000 204.320 2795.600 205.720 ;
        RECT 4.000 162.200 2796.000 204.320 ;
        RECT 4.000 160.800 2795.600 162.200 ;
        RECT 4.000 118.680 2796.000 160.800 ;
        RECT 4.000 117.280 2795.600 118.680 ;
        RECT 4.000 75.160 2796.000 117.280 ;
        RECT 4.000 73.760 2795.600 75.160 ;
        RECT 4.000 31.640 2796.000 73.760 ;
        RECT 4.000 30.240 2795.600 31.640 ;
        RECT 4.000 10.715 2796.000 30.240 ;
  END
END R4_butter
END LIBRARY

