magic
tech sky130A
magscale 1 2
timestamp 1699029394
<< obsli1 >>
rect 1104 2159 35236 36465
<< obsm1 >>
rect 474 892 35866 36496
<< metal2 >>
rect 478 0 534 800
rect 1214 0 1270 800
rect 1950 0 2006 800
rect 2686 0 2742 800
rect 3422 0 3478 800
rect 4158 0 4214 800
rect 4894 0 4950 800
rect 5630 0 5686 800
rect 6366 0 6422 800
rect 7102 0 7158 800
rect 7838 0 7894 800
rect 8574 0 8630 800
rect 9310 0 9366 800
rect 10046 0 10102 800
rect 10782 0 10838 800
rect 11518 0 11574 800
rect 12254 0 12310 800
rect 12990 0 13046 800
rect 13726 0 13782 800
rect 14462 0 14518 800
rect 15198 0 15254 800
rect 15934 0 15990 800
rect 16670 0 16726 800
rect 17406 0 17462 800
rect 18142 0 18198 800
rect 18878 0 18934 800
rect 19614 0 19670 800
rect 20350 0 20406 800
rect 21086 0 21142 800
rect 21822 0 21878 800
rect 22558 0 22614 800
rect 23294 0 23350 800
rect 24030 0 24086 800
rect 24766 0 24822 800
rect 25502 0 25558 800
rect 26238 0 26294 800
rect 26974 0 27030 800
rect 27710 0 27766 800
rect 28446 0 28502 800
rect 29182 0 29238 800
rect 29918 0 29974 800
rect 30654 0 30710 800
rect 31390 0 31446 800
rect 32126 0 32182 800
rect 32862 0 32918 800
rect 33598 0 33654 800
rect 34334 0 34390 800
rect 35070 0 35126 800
rect 35806 0 35862 800
<< obsm2 >>
rect 480 856 35860 36485
rect 590 734 1158 856
rect 1326 734 1894 856
rect 2062 734 2630 856
rect 2798 734 3366 856
rect 3534 734 4102 856
rect 4270 734 4838 856
rect 5006 734 5574 856
rect 5742 734 6310 856
rect 6478 734 7046 856
rect 7214 734 7782 856
rect 7950 734 8518 856
rect 8686 734 9254 856
rect 9422 734 9990 856
rect 10158 734 10726 856
rect 10894 734 11462 856
rect 11630 734 12198 856
rect 12366 734 12934 856
rect 13102 734 13670 856
rect 13838 734 14406 856
rect 14574 734 15142 856
rect 15310 734 15878 856
rect 16046 734 16614 856
rect 16782 734 17350 856
rect 17518 734 18086 856
rect 18254 734 18822 856
rect 18990 734 19558 856
rect 19726 734 20294 856
rect 20462 734 21030 856
rect 21198 734 21766 856
rect 21934 734 22502 856
rect 22670 734 23238 856
rect 23406 734 23974 856
rect 24142 734 24710 856
rect 24878 734 25446 856
rect 25614 734 26182 856
rect 26350 734 26918 856
rect 27086 734 27654 856
rect 27822 734 28390 856
rect 28558 734 29126 856
rect 29294 734 29862 856
rect 30030 734 30598 856
rect 30766 734 31334 856
rect 31502 734 32070 856
rect 32238 734 32806 856
rect 32974 734 33542 856
rect 33710 734 34278 856
rect 34446 734 35014 856
rect 35182 734 35750 856
<< metal3 >>
rect 35600 33736 36400 33856
rect 35600 24080 36400 24200
rect 35600 14424 36400 14544
rect 35600 4768 36400 4888
<< obsm3 >>
rect 4210 33936 35600 36481
rect 4210 33656 35520 33936
rect 4210 24280 35600 33656
rect 4210 24000 35520 24280
rect 4210 14624 35600 24000
rect 4210 14344 35520 14624
rect 4210 4968 35600 14344
rect 4210 4688 35520 4968
rect 4210 2143 35600 4688
<< metal4 >>
rect 4208 2128 4528 36496
rect 19568 2128 19888 36496
rect 34928 2128 35248 36496
<< labels >>
rlabel metal2 s 35806 0 35862 800 6 CLK
port 1 nsew signal input
rlabel metal3 s 35600 33736 36400 33856 6 RST
port 2 nsew signal input
rlabel metal2 s 24766 0 24822 800 6 Xio[0]
port 3 nsew signal output
rlabel metal2 s 26238 0 26294 800 6 Xio[1]
port 4 nsew signal output
rlabel metal2 s 27710 0 27766 800 6 Xio[2]
port 5 nsew signal output
rlabel metal2 s 29182 0 29238 800 6 Xio[3]
port 6 nsew signal output
rlabel metal2 s 24030 0 24086 800 6 Xro[0]
port 7 nsew signal output
rlabel metal2 s 25502 0 25558 800 6 Xro[1]
port 8 nsew signal output
rlabel metal2 s 26974 0 27030 800 6 Xro[2]
port 9 nsew signal output
rlabel metal2 s 28446 0 28502 800 6 Xro[3]
port 10 nsew signal output
rlabel metal3 s 35600 4768 36400 4888 6 c1
port 11 nsew signal input
rlabel metal3 s 35600 14424 36400 14544 6 c2
port 12 nsew signal input
rlabel metal3 s 35600 24080 36400 24200 6 c3
port 13 nsew signal input
rlabel metal2 s 29918 0 29974 800 6 la_oenb[0]
port 14 nsew signal output
rlabel metal2 s 30654 0 30710 800 6 la_oenb[1]
port 15 nsew signal output
rlabel metal2 s 31390 0 31446 800 6 la_oenb[2]
port 16 nsew signal output
rlabel metal2 s 32126 0 32182 800 6 la_oenb[3]
port 17 nsew signal output
rlabel metal2 s 32862 0 32918 800 6 la_oenb[4]
port 18 nsew signal output
rlabel metal2 s 33598 0 33654 800 6 la_oenb[5]
port 19 nsew signal output
rlabel metal2 s 34334 0 34390 800 6 la_oenb[6]
port 20 nsew signal output
rlabel metal2 s 35070 0 35126 800 6 la_oenb[7]
port 21 nsew signal output
rlabel metal4 s 4208 2128 4528 36496 6 vccd1
port 22 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 36496 6 vccd1
port 22 nsew power bidirectional
rlabel metal4 s 19568 2128 19888 36496 6 vssd1
port 23 nsew ground bidirectional
rlabel metal2 s 1214 0 1270 800 6 xi0[0]
port 24 nsew signal input
rlabel metal2 s 7102 0 7158 800 6 xi0[1]
port 25 nsew signal input
rlabel metal2 s 12990 0 13046 800 6 xi0[2]
port 26 nsew signal input
rlabel metal2 s 18878 0 18934 800 6 xi0[3]
port 27 nsew signal input
rlabel metal2 s 2686 0 2742 800 6 xi1[0]
port 28 nsew signal input
rlabel metal2 s 8574 0 8630 800 6 xi1[1]
port 29 nsew signal input
rlabel metal2 s 14462 0 14518 800 6 xi1[2]
port 30 nsew signal input
rlabel metal2 s 20350 0 20406 800 6 xi1[3]
port 31 nsew signal input
rlabel metal2 s 4158 0 4214 800 6 xi2[0]
port 32 nsew signal input
rlabel metal2 s 10046 0 10102 800 6 xi2[1]
port 33 nsew signal input
rlabel metal2 s 15934 0 15990 800 6 xi2[2]
port 34 nsew signal input
rlabel metal2 s 21822 0 21878 800 6 xi2[3]
port 35 nsew signal input
rlabel metal2 s 5630 0 5686 800 6 xi3[0]
port 36 nsew signal input
rlabel metal2 s 11518 0 11574 800 6 xi3[1]
port 37 nsew signal input
rlabel metal2 s 17406 0 17462 800 6 xi3[2]
port 38 nsew signal input
rlabel metal2 s 23294 0 23350 800 6 xi3[3]
port 39 nsew signal input
rlabel metal2 s 478 0 534 800 6 xr0[0]
port 40 nsew signal input
rlabel metal2 s 6366 0 6422 800 6 xr0[1]
port 41 nsew signal input
rlabel metal2 s 12254 0 12310 800 6 xr0[2]
port 42 nsew signal input
rlabel metal2 s 18142 0 18198 800 6 xr0[3]
port 43 nsew signal input
rlabel metal2 s 1950 0 2006 800 6 xr1[0]
port 44 nsew signal input
rlabel metal2 s 7838 0 7894 800 6 xr1[1]
port 45 nsew signal input
rlabel metal2 s 13726 0 13782 800 6 xr1[2]
port 46 nsew signal input
rlabel metal2 s 19614 0 19670 800 6 xr1[3]
port 47 nsew signal input
rlabel metal2 s 3422 0 3478 800 6 xr2[0]
port 48 nsew signal input
rlabel metal2 s 9310 0 9366 800 6 xr2[1]
port 49 nsew signal input
rlabel metal2 s 15198 0 15254 800 6 xr2[2]
port 50 nsew signal input
rlabel metal2 s 21086 0 21142 800 6 xr2[3]
port 51 nsew signal input
rlabel metal2 s 4894 0 4950 800 6 xr3[0]
port 52 nsew signal input
rlabel metal2 s 10782 0 10838 800 6 xr3[1]
port 53 nsew signal input
rlabel metal2 s 16670 0 16726 800 6 xr3[2]
port 54 nsew signal input
rlabel metal2 s 22558 0 22614 800 6 xr3[3]
port 55 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 36400 38800
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 509124
string GDS_FILE /home/guanyanlye/unic-cass/caravel_tutorial/caravel_user_example/openlane/R4_butter/runs/23_11_04_00_35/results/signoff/R4_butter.magic.gds
string GDS_START 79522
<< end >>

