magic
tech sky130A
magscale 1 2
timestamp 1696311228
<< obsli1 >>
rect 1104 2159 58880 37553
<< obsm1 >>
rect 934 2128 59050 37584
<< metal2 >>
rect 7470 0 7526 800
rect 22466 0 22522 800
rect 37462 0 37518 800
rect 52458 0 52514 800
<< obsm2 >>
rect 938 856 59046 38593
rect 938 800 7414 856
rect 7582 800 22410 856
rect 22578 800 37406 856
rect 37574 800 52402 856
rect 52570 800 59046 856
<< metal3 >>
rect 59200 38496 60000 38616
rect 59200 37544 60000 37664
rect 59200 36592 60000 36712
rect 59200 35640 60000 35760
rect 59200 34688 60000 34808
rect 59200 33736 60000 33856
rect 0 33192 800 33312
rect 59200 32784 60000 32904
rect 59200 31832 60000 31952
rect 59200 30880 60000 31000
rect 59200 29928 60000 30048
rect 59200 28976 60000 29096
rect 59200 28024 60000 28144
rect 59200 27072 60000 27192
rect 59200 26120 60000 26240
rect 59200 25168 60000 25288
rect 59200 24216 60000 24336
rect 59200 23264 60000 23384
rect 59200 22312 60000 22432
rect 59200 21360 60000 21480
rect 59200 20408 60000 20528
rect 0 19864 800 19984
rect 59200 19456 60000 19576
rect 59200 18504 60000 18624
rect 59200 17552 60000 17672
rect 59200 16600 60000 16720
rect 59200 15648 60000 15768
rect 59200 14696 60000 14816
rect 59200 13744 60000 13864
rect 59200 12792 60000 12912
rect 59200 11840 60000 11960
rect 59200 10888 60000 11008
rect 59200 9936 60000 10056
rect 59200 8984 60000 9104
rect 59200 8032 60000 8152
rect 59200 7080 60000 7200
rect 0 6536 800 6656
rect 59200 6128 60000 6248
rect 59200 5176 60000 5296
rect 59200 4224 60000 4344
rect 59200 3272 60000 3392
rect 59200 2320 60000 2440
rect 59200 1368 60000 1488
<< obsm3 >>
rect 800 38416 59120 38589
rect 800 37744 59200 38416
rect 800 37464 59120 37744
rect 800 36792 59200 37464
rect 800 36512 59120 36792
rect 800 35840 59200 36512
rect 800 35560 59120 35840
rect 800 34888 59200 35560
rect 800 34608 59120 34888
rect 800 33936 59200 34608
rect 800 33656 59120 33936
rect 800 33392 59200 33656
rect 880 33112 59200 33392
rect 800 32984 59200 33112
rect 800 32704 59120 32984
rect 800 32032 59200 32704
rect 800 31752 59120 32032
rect 800 31080 59200 31752
rect 800 30800 59120 31080
rect 800 30128 59200 30800
rect 800 29848 59120 30128
rect 800 29176 59200 29848
rect 800 28896 59120 29176
rect 800 28224 59200 28896
rect 800 27944 59120 28224
rect 800 27272 59200 27944
rect 800 26992 59120 27272
rect 800 26320 59200 26992
rect 800 26040 59120 26320
rect 800 25368 59200 26040
rect 800 25088 59120 25368
rect 800 24416 59200 25088
rect 800 24136 59120 24416
rect 800 23464 59200 24136
rect 800 23184 59120 23464
rect 800 22512 59200 23184
rect 800 22232 59120 22512
rect 800 21560 59200 22232
rect 800 21280 59120 21560
rect 800 20608 59200 21280
rect 800 20328 59120 20608
rect 800 20064 59200 20328
rect 880 19784 59200 20064
rect 800 19656 59200 19784
rect 800 19376 59120 19656
rect 800 18704 59200 19376
rect 800 18424 59120 18704
rect 800 17752 59200 18424
rect 800 17472 59120 17752
rect 800 16800 59200 17472
rect 800 16520 59120 16800
rect 800 15848 59200 16520
rect 800 15568 59120 15848
rect 800 14896 59200 15568
rect 800 14616 59120 14896
rect 800 13944 59200 14616
rect 800 13664 59120 13944
rect 800 12992 59200 13664
rect 800 12712 59120 12992
rect 800 12040 59200 12712
rect 800 11760 59120 12040
rect 800 11088 59200 11760
rect 800 10808 59120 11088
rect 800 10136 59200 10808
rect 800 9856 59120 10136
rect 800 9184 59200 9856
rect 800 8904 59120 9184
rect 800 8232 59200 8904
rect 800 7952 59120 8232
rect 800 7280 59200 7952
rect 800 7000 59120 7280
rect 800 6736 59200 7000
rect 880 6456 59200 6736
rect 800 6328 59200 6456
rect 800 6048 59120 6328
rect 800 5376 59200 6048
rect 800 5096 59120 5376
rect 800 4424 59200 5096
rect 800 4144 59120 4424
rect 800 3472 59200 4144
rect 800 3192 59120 3472
rect 800 2520 59200 3192
rect 800 2240 59120 2520
rect 800 1568 59200 2240
rect 800 1395 59120 1568
<< metal4 >>
rect 4208 2128 4528 37584
rect 19568 2128 19888 37584
rect 34928 2128 35248 37584
rect 50288 2128 50608 37584
<< labels >>
rlabel metal3 s 59200 9936 60000 10056 6 Xio[0]
port 1 nsew signal output
rlabel metal3 s 59200 19456 60000 19576 6 Xio[1]
port 2 nsew signal output
rlabel metal3 s 59200 28976 60000 29096 6 Xio[2]
port 3 nsew signal output
rlabel metal3 s 59200 38496 60000 38616 6 Xio[3]
port 4 nsew signal output
rlabel metal3 s 59200 8984 60000 9104 6 Xro[0]
port 5 nsew signal output
rlabel metal3 s 59200 18504 60000 18624 6 Xro[1]
port 6 nsew signal output
rlabel metal3 s 59200 28024 60000 28144 6 Xro[2]
port 7 nsew signal output
rlabel metal3 s 59200 37544 60000 37664 6 Xro[3]
port 8 nsew signal output
rlabel metal3 s 0 33192 800 33312 6 c1
port 9 nsew signal input
rlabel metal3 s 0 19864 800 19984 6 c2
port 10 nsew signal input
rlabel metal3 s 0 6536 800 6656 6 c3
port 11 nsew signal input
rlabel metal2 s 7470 0 7526 800 6 la_oenb[0]
port 12 nsew signal output
rlabel metal2 s 22466 0 22522 800 6 la_oenb[1]
port 13 nsew signal output
rlabel metal2 s 37462 0 37518 800 6 la_oenb[2]
port 14 nsew signal output
rlabel metal2 s 52458 0 52514 800 6 la_oenb[3]
port 15 nsew signal output
rlabel metal4 s 4208 2128 4528 37584 6 vccd1
port 16 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 37584 6 vccd1
port 16 nsew power bidirectional
rlabel metal4 s 19568 2128 19888 37584 6 vssd1
port 17 nsew ground bidirectional
rlabel metal4 s 50288 2128 50608 37584 6 vssd1
port 17 nsew ground bidirectional
rlabel metal3 s 59200 2320 60000 2440 6 xi0[0]
port 18 nsew signal input
rlabel metal3 s 59200 11840 60000 11960 6 xi0[1]
port 19 nsew signal input
rlabel metal3 s 59200 21360 60000 21480 6 xi0[2]
port 20 nsew signal input
rlabel metal3 s 59200 30880 60000 31000 6 xi0[3]
port 21 nsew signal input
rlabel metal3 s 59200 4224 60000 4344 6 xi1[0]
port 22 nsew signal input
rlabel metal3 s 59200 13744 60000 13864 6 xi1[1]
port 23 nsew signal input
rlabel metal3 s 59200 23264 60000 23384 6 xi1[2]
port 24 nsew signal input
rlabel metal3 s 59200 32784 60000 32904 6 xi1[3]
port 25 nsew signal input
rlabel metal3 s 59200 6128 60000 6248 6 xi2[0]
port 26 nsew signal input
rlabel metal3 s 59200 15648 60000 15768 6 xi2[1]
port 27 nsew signal input
rlabel metal3 s 59200 25168 60000 25288 6 xi2[2]
port 28 nsew signal input
rlabel metal3 s 59200 34688 60000 34808 6 xi2[3]
port 29 nsew signal input
rlabel metal3 s 59200 8032 60000 8152 6 xi3[0]
port 30 nsew signal input
rlabel metal3 s 59200 17552 60000 17672 6 xi3[1]
port 31 nsew signal input
rlabel metal3 s 59200 27072 60000 27192 6 xi3[2]
port 32 nsew signal input
rlabel metal3 s 59200 36592 60000 36712 6 xi3[3]
port 33 nsew signal input
rlabel metal3 s 59200 1368 60000 1488 6 xr0[0]
port 34 nsew signal input
rlabel metal3 s 59200 10888 60000 11008 6 xr0[1]
port 35 nsew signal input
rlabel metal3 s 59200 20408 60000 20528 6 xr0[2]
port 36 nsew signal input
rlabel metal3 s 59200 29928 60000 30048 6 xr0[3]
port 37 nsew signal input
rlabel metal3 s 59200 3272 60000 3392 6 xr1[0]
port 38 nsew signal input
rlabel metal3 s 59200 12792 60000 12912 6 xr1[1]
port 39 nsew signal input
rlabel metal3 s 59200 22312 60000 22432 6 xr1[2]
port 40 nsew signal input
rlabel metal3 s 59200 31832 60000 31952 6 xr1[3]
port 41 nsew signal input
rlabel metal3 s 59200 5176 60000 5296 6 xr2[0]
port 42 nsew signal input
rlabel metal3 s 59200 14696 60000 14816 6 xr2[1]
port 43 nsew signal input
rlabel metal3 s 59200 24216 60000 24336 6 xr2[2]
port 44 nsew signal input
rlabel metal3 s 59200 33736 60000 33856 6 xr2[3]
port 45 nsew signal input
rlabel metal3 s 59200 7080 60000 7200 6 xr3[0]
port 46 nsew signal input
rlabel metal3 s 59200 16600 60000 16720 6 xr3[1]
port 47 nsew signal input
rlabel metal3 s 59200 26120 60000 26240 6 xr3[2]
port 48 nsew signal input
rlabel metal3 s 59200 35640 60000 35760 6 xr3[3]
port 49 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 60000 40000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 645856
string GDS_FILE /home/guanyanlye/unic-cass/caravel_tutorial/caravel_uniccas_example/openlane/R4_butter/runs/23_10_03_13_32/results/signoff/R4_butter.magic.gds
string GDS_START 53070
<< end >>

